module leading_one_div(
input [23:0] A,
output [4:0] msb_loc
);

assign msb_loc = (A[23]==1) ? 23 : (A[22]==1) ? 22 : (A[21]==1) ? 21 : (A[20]==1) ? 20 : (A[19]==1) ? 19 : (A[18]==1) ? 18 : (A[17]==1) ? 17 : (A[16]==1) ? 16 : (A[15]==1) ? 15 : (A[14]==1) ? 14 : (A[13]==1) ? 13 : (A[12]==1) ? 12 : (A[11]==1) ? 11 : (A[10]==1) ? 10 : (A[9]==1) ? 9 : (A[8]==1) ? 8 : (A[7]==1) ? 7 : (A[6]==1) ? 6 : (A[5]==1) ? 5 : (A[4]==1) ? 4 : (A[3]==1) ? 3 : (A[2]==1) ? 2 : (A[1]==1) ? 1 : 0;

endmodule
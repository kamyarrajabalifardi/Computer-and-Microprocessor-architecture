module leading_one(
input [48:0] A,
output [5:0] msb_loc
);

assign msb_loc = (A[48] == 1) ? 48 : (A[47]==1) ? 47 : (A[46]==1) ? 46 : (A[45]==1) ? 45 : (A[44]==1) ? 44 : (A[43]==1) ? 43 : (A[42]==1) ? 42 : (A[41]==1) ? 41 : (A[40]==1) ? 40 : (A[39]==1) ? 39 : (A[38]==1) ? 38 : (A[37]==1) ? 37 : (A[36]==1) ? 36 : (A[35]==1) ? 35 : (A[34]==1) ? 34 : (A[33]==1) ? 33 : (A[32]==1) ? 32 : (A[31]==1) ? 31 : (A[30]==1) ? 30 : (A[29]==1) ? 29 : (A[28]==1) ? 28 : (A[28]==1) ? 28 : (A[27]==1) ? 27 : (A[26]==1) ? 26 : (A[25]==1) ? 25 : (A[24]==1) ? 24 : (A[23]==1) ? 23 : (A[22]==1) ? 22 : (A[21]==1) ? 21 : (A[20]==1) ? 20 : (A[19]==1) ? 19 : (A[18]==1) ? 18 : (A[17]==1) ? 17 : (A[16]==1) ? 16 : (A[15]==1) ? 15 : (A[14]==1) ? 14 : (A[13]==1) ? 13 : (A[12]==1) ? 12 : (A[11]==1) ? 11 : (A[10]==1) ? 10 : (A[9]==1) ? 9 : (A[8]==1) ? 8 : (A[7]==1) ? 7 : (A[6]==1) ? 6 : (A[5]==1) ? 5 : (A[4]==1) ? 4 : (A[3]==1) ? 3 : (A[2]==1) ? 2 : (A[1]==1) ? 1 : 0;

endmodule